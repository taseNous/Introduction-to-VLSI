CIRCUIT D:\Documents and Settings\sicard\Mes documents\microwind31\examples\InvCapa.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
Vin 5 0 DC 0 PULSE(0.00 1.20 0.98N 0.02N 0.02N 0.98N 2.00N)
*
* List of nodes
* "inv" corresponds to n�3
* "in" corresponds to n�5
*
* MOS devices
MN1 0 5 3 0 N1  W= 0.24U L= 0.12U
MP1 1 5 3 1 P1  W= 0.24U L= 0.12U
*
C2 1 0  1.256fF
C3 3 0  0.487fF
C5 5 0  0.314fF
*
* Extra RLC
*
Cadd1 3 0 0.01pF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTHO=0.40 U0=0.050 TOXE= 2.0E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.050 UA=3.000e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTHO=-0.45 U0=0.018 TOXE= 2.0E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.018 UA=1.500e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p
*
* Transient analysis
*
* (Winspice)
.options temp=27.0
.control
tran 0.1N 5.00N
print  V(5) V(3) > out.txt
plot  V(5) V(3)
.endc
.END
